module top_module (MAX10_CLK1_50, KEY, HEX0, HEX1, HEX2, HEX3,LEDR);
input [1:0] KEY;
input MAX10_CLK1_50;
output [6:0] HEX0, HEX1, HEX2, HEX3;
output [9:0] LEDR;

endmodule //top_module
