module top_module ();

endmodule //
