module BCD_counter ();

endmodule //BCD_counter
