module BCD_decoder ();
4'b0000:HEXx[6:0] = 7'b1000000;
4'b0001:HEXx[6:0] = 7'b1111001;
4'b0010:HEXx[6:0] = 7'b0100100;
4'b0011:HEXx[6:0] = 7'b0110000;
4'b0100:HEXx[6:0] = 7'b0011001;
4'b0101:HEXx[6:0] = 7'b0010010;
4'b0110:HEXx[6:0] = 7'b0000010;
4'b0111:HEXx[6:0] = 7'b1111000;
4'b1000:HEXx[6:0] = 7'b0000000;
4'b1001:HEXx[6:0] = 7'b0011000;
endmodule //BCD_decoder
