module BCD_decoder ();

endmodule //BCD_decoder
