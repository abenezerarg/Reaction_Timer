module Clock_divider ();

endmodule //Clock_divider
