module LFSR ();

endmodule //LFSR
